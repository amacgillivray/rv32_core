`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: EECS 581 Team 11
// Engineer: Andrew MacGillivray
// 
// Create Date: 11/20/2022 03:37:49 PM
// Design Name: CSR Unit
// Module Name: csr
// Project Name: Linear Algebra Accelerator
// Target Devices: 
// Description: 
// 
// Revision:
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module csr(
    input [31:0] pc
);
    reg[31:0] scause;
    reg[31:0] sepc;
    // todo: behavior
endmodule