`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: EECS 581 Team 11
// Engineer: Jarrod Grothusen
// 
// Create Date: 
// Design Name: 
// Module Name: ex_ALU_frwd
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ex_ALU_frwd(
    input ctrl_mux4,
    input ctrl_mux3,
    input idex_regRS1,
    input idex_regRS2,
    output exmem_regRD,
    output exmem_regWrite,
    output memwb_regRD,
    output memwb_regWrite
    );
    
endmodule
