`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: EECS 581 Team 11
// Engineer: Andrew MacGillivray
// 
// Create Date: 10/29/2022 01:13:53 PM
// Design Name: 
// Module Name: forwarding_unit_branch
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module forwarding_unit_branch(
    output ctrl_mux_1_branch,
    output ctrl_mux_2_branch,
    input IFID_Reg_RS1,
    input IFID_Reg_RS2,
    input EXMEM_Reg_RD,
    input EXMEM_MemToReg
    );
endmodule
